-- Testbench float16 random pseudonym without NaN/Inf/overflow/underflow
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

constant NUM_CYCLES : integer := 16;
type float_array is array (0 to NUM_CYCLES-1) of std_logic_vector(15 downto 0);

constant input_A : float_array := (
    "1010110010111101",
    "0100100011011011",
    "0100001110000111",
    "0100011010111000",
    "1100010000000101",
    "1011100010001011",
    "0100010100110110",
    "0100100001010000",
    "0100000110001100",
    "1010110111000101",
    "1100100000110001",
    "0100010100001101",
    "0100010010011010",
    "0011010000100111",
    "0100001111110000",
    "0011110011000001"
);

constant input_B : float_array := (
    "1100011010010111",
    "0100100010010001",
    "0100100001000101",
    "0100000101000000",
    "0011111011010101",
    "1100001001000001",
    "1100010101001010",
    "1100000111111100",
    "0100000101010101",
    "1100011100111111",
    "1100011011001011",
    "1100100010010111",
    "1100100001101110",
    "0100001010001000",
    "0100000110101010",
    "1011100101101010"
);

constant expected_result : std_logic_vector(15 downto 0) := "0101010001011010";
